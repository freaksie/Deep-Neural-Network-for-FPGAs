reg [(10-1):0] ram [0:(1024-1)] = '{10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h000
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h001
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h002
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h003
,10'h004
,10'h004
,10'h004
,10'h004
,10'h004
,10'h004
,10'h004
,10'h004
,10'h004
,10'h004
,10'h004
,10'h004
,10'h004
,10'h004
,10'h005
,10'h005
,10'h005
,10'h005
,10'h005
,10'h005
,10'h005
,10'h005
,10'h005
,10'h005
,10'h005
,10'h005
,10'h006
,10'h006
,10'h006
,10'h006
,10'h006
,10'h006
,10'h006
,10'h006
,10'h006
,10'h006
,10'h007
,10'h007
,10'h007
,10'h007
,10'h007
,10'h007
,10'h007
,10'h007
,10'h008
,10'h008
,10'h008
,10'h008
,10'h008
,10'h008
,10'h008
,10'h008
,10'h009
,10'h009
,10'h009
,10'h009
,10'h009
,10'h009
,10'h009
,10'h00A
,10'h00A
,10'h00A
,10'h00A
,10'h00A
,10'h00A
,10'h00B
,10'h00B
,10'h00B
,10'h00B
,10'h00B
,10'h00B
,10'h00C
,10'h00C
,10'h00C
,10'h00C
,10'h00C
,10'h00D
,10'h00D
,10'h00D
,10'h00D
,10'h00D
,10'h00E
,10'h00E
,10'h00E
,10'h00E
,10'h00F
,10'h00F
,10'h00F
,10'h00F
,10'h010
,10'h010
,10'h010
,10'h010
,10'h011
,10'h011
,10'h011
,10'h011
,10'h012
,10'h012
,10'h012
,10'h012
,10'h013
,10'h013
,10'h013
,10'h014
,10'h014
,10'h014
,10'h015
,10'h015
,10'h015
,10'h016
,10'h016
,10'h016
,10'h017
,10'h017
,10'h017
,10'h018
,10'h018
,10'h019
,10'h019
,10'h019
,10'h01A
,10'h01A
,10'h01A
,10'h01B
,10'h01B
,10'h01C
,10'h01C
,10'h01D
,10'h01D
,10'h01E
,10'h01E
,10'h01E
,10'h01F
,10'h01F
,10'h020
,10'h020
,10'h021
,10'h021
,10'h022
,10'h022
,10'h023
,10'h023
,10'h024
,10'h025
,10'h025
,10'h026
,10'h026
,10'h027
,10'h027
,10'h028
,10'h029
,10'h029
,10'h02A
,10'h02B
,10'h02B
,10'h02C
,10'h02D
,10'h02D
,10'h02E
,10'h02F
,10'h02F
,10'h030
,10'h031
,10'h032
,10'h032
,10'h033
,10'h034
,10'h035
,10'h035
,10'h036
,10'h037
,10'h038
,10'h039
,10'h03A
,10'h03A
,10'h03B
,10'h03C
,10'h03D
,10'h03E
,10'h03F
,10'h040
,10'h041
,10'h042
,10'h043
,10'h044
,10'h045
,10'h046
,10'h047
,10'h048
,10'h049
,10'h04A
,10'h04B
,10'h04C
,10'h04D
,10'h04E
,10'h04F
,10'h051
,10'h052
,10'h053
,10'h054
,10'h055
,10'h057
,10'h058
,10'h059
,10'h05A
,10'h05C
,10'h05D
,10'h05E
,10'h060
,10'h061
,10'h063
,10'h064
,10'h065
,10'h067
,10'h068
,10'h06A
,10'h06B
,10'h06D
,10'h06E
,10'h070
,10'h071
,10'h073
,10'h075
,10'h076
,10'h078
,10'h07A
,10'h07B
,10'h07D
,10'h07F
,10'h080
,10'h082
,10'h084
,10'h086
,10'h088
,10'h08A
,10'h08B
,10'h08D
,10'h08F
,10'h091
,10'h093
,10'h095
,10'h097
,10'h099
,10'h09B
,10'h09D
,10'h09F
,10'h0A1
,10'h0A4
,10'h0A6
,10'h0A8
,10'h0AA
,10'h0AC
,10'h0AF
,10'h0B1
,10'h0B3
,10'h0B6
,10'h0B8
,10'h0BA
,10'h0BD
,10'h0BF
,10'h0C2
,10'h0C4
,10'h0C7
,10'h0C9
,10'h0CC
,10'h0CE
,10'h0D1
,10'h0D3
,10'h0D6
,10'h0D9
,10'h0DB
,10'h0DE
,10'h0E1
,10'h0E4
,10'h0E6
,10'h0E9
,10'h0EC
,10'h0EF
,10'h0F2
,10'h0F5
,10'h0F8
,10'h0FA
,10'h0FD
,10'h100
,10'h103
,10'h106
,10'h10A
,10'h10D
,10'h110
,10'h113
,10'h116
,10'h119
,10'h11C
,10'h120
,10'h123
,10'h126
,10'h129
,10'h12D
,10'h130
,10'h133
,10'h137
,10'h13A
,10'h13E
,10'h141
,10'h145
,10'h148
,10'h14C
,10'h14F
,10'h153
,10'h156
,10'h15A
,10'h15D
,10'h161
,10'h165
,10'h168
,10'h16C
,10'h16F
,10'h173
,10'h177
,10'h17B
,10'h17E
,10'h182
,10'h186
,10'h18A
,10'h18D
,10'h191
,10'h195
,10'h199
,10'h19D
,10'h1A1
,10'h1A4
,10'h1A8
,10'h1AC
,10'h1B0
,10'h1B4
,10'h1B8
,10'h1BC
,10'h1C0
,10'h1C4
,10'h1C8
,10'h1CC
,10'h1D0
,10'h1D4
,10'h1D8
,10'h1DC
,10'h1E0
,10'h1E4
,10'h1E8
,10'h1EC
,10'h1F0
,10'h1F4
,10'h1F8
,10'h1FC
,10'h200
,10'h203
,10'h207
,10'h20B
,10'h20F
,10'h213
,10'h217
,10'h21B
,10'h21F
,10'h223
,10'h227
,10'h22B
,10'h22F
,10'h233
,10'h237
,10'h23B
,10'h23F
,10'h243
,10'h247
,10'h24B
,10'h24F
,10'h253
,10'h257
,10'h25B
,10'h25E
,10'h262
,10'h266
,10'h26A
,10'h26E
,10'h272
,10'h275
,10'h279
,10'h27D
,10'h281
,10'h284
,10'h288
,10'h28C
,10'h290
,10'h293
,10'h297
,10'h29A
,10'h29E
,10'h2A2
,10'h2A5
,10'h2A9
,10'h2AC
,10'h2B0
,10'h2B3
,10'h2B7
,10'h2BA
,10'h2BE
,10'h2C1
,10'h2C5
,10'h2C8
,10'h2CC
,10'h2CF
,10'h2D2
,10'h2D6
,10'h2D9
,10'h2DC
,10'h2DF
,10'h2E3
,10'h2E6
,10'h2E9
,10'h2EC
,10'h2EF
,10'h2F2
,10'h2F5
,10'h2F9
,10'h2FC
,10'h2FF
,10'h302
,10'h305
,10'h307
,10'h30A
,10'h30D
,10'h310
,10'h313
,10'h316
,10'h319
,10'h31B
,10'h31E
,10'h321
,10'h324
,10'h326
,10'h329
,10'h32C
,10'h32E
,10'h331
,10'h333
,10'h336
,10'h338
,10'h33B
,10'h33D
,10'h340
,10'h342
,10'h345
,10'h347
,10'h349
,10'h34C
,10'h34E
,10'h350
,10'h353
,10'h355
,10'h357
,10'h359
,10'h35B
,10'h35E
,10'h360
,10'h362
,10'h364
,10'h366
,10'h368
,10'h36A
,10'h36C
,10'h36E
,10'h370
,10'h372
,10'h374
,10'h375
,10'h377
,10'h379
,10'h37B
,10'h37D
,10'h37F
,10'h380
,10'h382
,10'h384
,10'h385
,10'h387
,10'h389
,10'h38A
,10'h38C
,10'h38E
,10'h38F
,10'h391
,10'h392
,10'h394
,10'h395
,10'h397
,10'h398
,10'h39A
,10'h39B
,10'h39C
,10'h39E
,10'h39F
,10'h3A1
,10'h3A2
,10'h3A3
,10'h3A5
,10'h3A6
,10'h3A7
,10'h3A8
,10'h3AA
,10'h3AB
,10'h3AC
,10'h3AD
,10'h3AE
,10'h3B0
,10'h3B1
,10'h3B2
,10'h3B3
,10'h3B4
,10'h3B5
,10'h3B6
,10'h3B7
,10'h3B8
,10'h3B9
,10'h3BA
,10'h3BB
,10'h3BC
,10'h3BD
,10'h3BE
,10'h3BF
,10'h3C0
,10'h3C1
,10'h3C2
,10'h3C3
,10'h3C4
,10'h3C5
,10'h3C5
,10'h3C6
,10'h3C7
,10'h3C8
,10'h3C9
,10'h3CA
,10'h3CA
,10'h3CB
,10'h3CC
,10'h3CD
,10'h3CD
,10'h3CE
,10'h3CF
,10'h3D0
,10'h3D0
,10'h3D1
,10'h3D2
,10'h3D2
,10'h3D3
,10'h3D4
,10'h3D4
,10'h3D5
,10'h3D6
,10'h3D6
,10'h3D7
,10'h3D8
,10'h3D8
,10'h3D9
,10'h3D9
,10'h3DA
,10'h3DA
,10'h3DB
,10'h3DC
,10'h3DC
,10'h3DD
,10'h3DD
,10'h3DE
,10'h3DE
,10'h3DF
,10'h3DF
,10'h3E0
,10'h3E0
,10'h3E1
,10'h3E1
,10'h3E1
,10'h3E2
,10'h3E2
,10'h3E3
,10'h3E3
,10'h3E4
,10'h3E4
,10'h3E5
,10'h3E5
,10'h3E5
,10'h3E6
,10'h3E6
,10'h3E6
,10'h3E7
,10'h3E7
,10'h3E8
,10'h3E8
,10'h3E8
,10'h3E9
,10'h3E9
,10'h3E9
,10'h3EA
,10'h3EA
,10'h3EA
,10'h3EB
,10'h3EB
,10'h3EB
,10'h3EC
,10'h3EC
,10'h3EC
,10'h3ED
,10'h3ED
,10'h3ED
,10'h3ED
,10'h3EE
,10'h3EE
,10'h3EE
,10'h3EE
,10'h3EF
,10'h3EF
,10'h3EF
,10'h3EF
,10'h3F0
,10'h3F0
,10'h3F0
,10'h3F0
,10'h3F1
,10'h3F1
,10'h3F1
,10'h3F1
,10'h3F2
,10'h3F2
,10'h3F2
,10'h3F2
,10'h3F2
,10'h3F3
,10'h3F3
,10'h3F3
,10'h3F3
,10'h3F3
,10'h3F4
,10'h3F4
,10'h3F4
,10'h3F4
,10'h3F4
,10'h3F4
,10'h3F5
,10'h3F5
,10'h3F5
,10'h3F5
,10'h3F5
,10'h3F5
,10'h3F6
,10'h3F6
,10'h3F6
,10'h3F6
,10'h3F6
,10'h3F6
,10'h3F6
,10'h3F7
,10'h3F7
,10'h3F7
,10'h3F7
,10'h3F7
,10'h3F7
,10'h3F7
,10'h3F7
,10'h3F8
,10'h3F8
,10'h3F8
,10'h3F8
,10'h3F8
,10'h3F8
,10'h3F8
,10'h3F8
,10'h3F9
,10'h3F9
,10'h3F9
,10'h3F9
,10'h3F9
,10'h3F9
,10'h3F9
,10'h3F9
,10'h3F9
,10'h3F9
,10'h3FA
,10'h3FA
,10'h3FA
,10'h3FA
,10'h3FA
,10'h3FA
,10'h3FA
,10'h3FA
,10'h3FA
,10'h3FA
,10'h3FA
,10'h3FA
,10'h3FB
,10'h3FB
,10'h3FB
,10'h3FB
,10'h3FB
,10'h3FB
,10'h3FB
,10'h3FB
,10'h3FB
,10'h3FB
,10'h3FB
,10'h3FB
,10'h3FB
,10'h3FB
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FC
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FD
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FE
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
,10'h3FF
};
